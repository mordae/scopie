*****************************************************
* Collection of SPICE models for the SinPI project *
*****************************************************
*
* Most models were written in 2022 by Jan Hamal Dvořák <mordae@anilinux.org>.
* Universal Op-Amp was written in 2019 by Ste Kulov, HD Retrovision LLC.
*
* To the extent possible under law, the author(s) have dedicated all copyright
* and related and neighboring rights to this software to the public domain worldwide.
* This software is distributed without any warranty.
* You should have received a copy of the CC0 Public Domain Dedication along with this software.
* If not, see <http://creativecommons.org/publicdomain/zero/1.0/>.
*

******************************************************************************
* Ideal gate that open at 1.2V with 0.8V hysteresis
******************************************************************************

.subckt IDEAL_GATE in out v+ v-
Sgate in out v+ v- gate ON
.model gate sw(vt=1.2, vh=0.8, ron=1u, roff=1G)
.ends


******************************************************************************
* Ideal AND gate with 50k pull-down
******************************************************************************

.subckt IDEAL_AND left right out v+ v-
X1 v+ tmp1 left v- IDEAL_GATE
X2 tmp1 out right v- IDEAL_GATE
R1 v- out 50k
.ends


******************************************************************************
* Ideal NOT gate with 50k pull-up
******************************************************************************

.subckt IDEAL_NOT in out v+ v-
X1 v- out in v- IDEAL_GATE
R1 v+ out 50k
.ends


******************************************************************************
* Ideal OR gate with 50k pull-up
******************************************************************************

.subckt IDEAL_OR left right out v+ v-
X1 left tmp v+ v- IDEAL_NOT
X2 right tmp v+ v- IDEAL_NOT
X3 tmp out v+ v- IDEAL_NOT
.ends


******************************************************************************
* 2P4T analog multiplexer
* Ideal model without delays
******************************************************************************

.subckt DG4052EEN-T1-GE4 y y3 y1 en v- gnd b a x3 x0 x x1 x2 v+ y0 y2
Rx rx x 80
Ry ry y 80

Cx gnd x 10p
Cy gnd y 10p

Cx0 gnd x0 2p
Cx1 gnd x0 2p
Cx2 gnd x0 2p
Cx3 gnd x0 2p

Cy0 gnd y0 2p
Cy1 gnd y0 2p
Cy2 gnd y0 2p
Cy3 gnd y0 2p

Xx0 x0 rx code0 gnd IDEAL_GATE
Xy0 y0 ry code0 gnd IDEAL_GATE

Xx1 x1 rx code1 gnd IDEAL_GATE
Xy1 y1 ry code1 gnd IDEAL_GATE

Xx2 x2 rx code2 gnd IDEAL_GATE
Xy2 y2 ry code2 gnd IDEAL_GATE

Xx3 x3 rx code3 gnd IDEAL_GATE
Xy3 y3 ry code3 gnd IDEAL_GATE

Xnota ra nota v+ v- IDEAL_NOT
Xnotb rb notb v+ v- IDEAL_NOT

Xcode0 nota notb code0 v+ gnd IDEAL_AND
Xcode1 nota   rb code1 v+ gnd IDEAL_AND
Xcode2   ra notb code2 v+ gnd IDEAL_AND
Xcode3   ra   rb code3 v+ gnd IDEAL_AND

Ra ra a 200k
Ca ra gnd 3.4p

Rb rb b 200k
Cb rb gnd 3.4p

* 1mA @ 10MHz v+ to v- @ 10V
Rp1 v+ v- 10k

* 100uA @ 10MHz v+ / v- to gnd @ 10V
Rp2 v+ gnd 100k
Rp3 v- gnd 100k

* enable pin pulls up the switches
Ren0 en code0 200k
Ren1 en code1 200k
Ren2 en code2 200k
Ren3 en code3 200k
.ends


******************************************************************************
* Two channel opamp with variable attenuator
******************************************************************************

.subckt LMH6521 A3 A4 A5 MOD0 MOD1 B5 B4 B3 B2 B1 INB+ INB- GND V+ GND B0 OUTB+ OUTB- ENB LATB LATA ENA OUTA- OUTA+ A0 GND V+ GND INA- INA+ A1 A2 GND
.param ata = 0
.param atb = 0

* Pull-ups on the unimportant pins we do not simulate.
Rlata LATA V+ 50k
Rlatb LATB V+ 50k
Rmod0 MOD0 V+ 50k
Rmod1 MOD1 V+ 50k
Ra0 A0 V+ 50k
Ra1 A1 V+ 50k
Ra2 A2 V+ 50k
Ra3 A3 V+ 50k
Ra4 A4 V+ 50k
Ra5 A5 V+ 50k
Rb0 B0 V+ 50k
Rb1 B1 V+ 50k
Rb2 B2 V+ 50k
Rb3 B3 V+ 50k
Rb4 B4 V+ 50k
Rb5 B5 V+ 50k
Rena ENA V+ 50k
Renb ENB V+ 50k

XA OUTA+ OUTA- INA+ INA- V+ GND LMH6521_CH at={ata}
XB OUTB+ OUTB- INB+ INB- V+ GND LMH6521_CH at={atb}
.ends LMH6521


* Single channel of the LMH6521 dual opamp
.subckt LMH6521_CH out+ out- in+ in- v+ gnd
.param at = 0

* Input resistances
Rrin+ in+ rin+ 200
Rrin- in- rin- 200

* Output resistances
Rrout+ out+ rout+ 20
Rrout- out- rout- 20

* Slight input bias
Rbias+v rin+ v+ 1Meg
Rbias+g rin+ gnd 1Meg
Rbias-v rin- v+ 1Meg
Rbias-g rin- gnd 1Meg

* Wing some parasitics
CPrin+ in+ gnd 1p
CPrin- in- gnd 1p
CProut+ out+ gnd 1p
CProut- out- gnd 1p

* Attenuator / Amplifier
Eamp rout+ rout- rin+ rin- {pwr(10, -at / 20) * pwr(10, 26 / 20)}

* Input voltage clamps
Din+1 rin+ v+ diode
Din+2 gnd rin+ diode
Din-1 rin- v+ diode
Din-2 gnd rin- diode

* Output voltage clamps
Dout+1 rout+ v+ diode
Dout+2 gnd out+ diode
Dout-1 rout- v+ diode
Dout-2 gnd out- diode

.model diode D(Is=1e-14)
.ends LMH6521_CH


******************************************************************************
*
* Universal Op-Amp
* Single pole opamp with rail saturation, current consumption,
* current limiting, and input offset voltage
*
* PINOUT ORDER  1   2   3   4   5
* PINOUT ORDER +IN -IN OUT VCC VEE
*
* Parameters:
* Avol => open-loop voltage gain (V/V), default=100k
* GBW => gain-bandwidth product (Hz), default=100meg
* Rin => differential input resistance (ohm), default=100g
* Rout => open-loop output resistance (ohm), default=1
* Iq => quiescent supply current (A), default=1m
* Ilimit => maximum output current (A), default=1
* Vrail => voltage between output saturation and each rail (V), default=0
* Vos => input offset voltage (V), default=0
* Vmax => total maximum supply voltage between rails (V), default=50
*
******************************************************************************

.subckt UOPAMP in+ in- out v+ v-
.param Avol=100k
.param GBW=100meg
.param Rin = 100g
.param Rout = 1
.param Iq = 1m
.param Ilimit = 1
.param Vrail = 0
.param Vos = 0
.param Vmax = 50
.param PI = 3.1415926535898
G1 v+ n1 offset in- 1u
G2 v- n1 offset in- 1u
R1 v+ n1 {Avol/1u}
R2 n1 v- {Avol/1u}
G3 out v+ v+ n1 {1/(2*Rout)}
G4 v- out n1 v- {1/(2*Rout)}
R4 v+ out {2*Rout}
R5 out v- {2*Rout}
C1 v+ n1 {1u/(2*PI*GBW)}
C2 n1 v- {1u/(2*PI*GBW)}
G6 n5 v- n1 out {1/(2*Rout)}
G5 n6 v- out n1 {1/(2*Rout)}
R8 in- in+ {Rin}
Vclamp+ v+ clamp+ {Vrail+545m}
Vclamp- clamp- v- {Vrail+545m}
Voffset offset in+ {Vos}
Vlimit- out limit- {Ilimit-545m}
Vlimit+ limit+ out {Ilimit-545m}
D1 n1 clamp+ diode
D2 clamp- n1 diode
D3 v+ n5 diode
D4 v+ n6 diode
D5 v- n5 zener
D6 v- n6 zener
D7 n1 limit+ diode
D8 limit- n1 diode
I1 v+ v- {Iq}
.model diode D(Is=1e-14)
.model zener D(Is=1e-14 BV={Vmax})
.ends


******************************************************************************
* Rectifier Diode
******************************************************************************

.subckt RRE04EA6DFH a1 nc a2 c1 c2
D1 a1 c1 diode
D2 a2 c2 diode
C1 a1 c1 1.2p
C2 a2 c2 1.2p
.model diode D(BV=600)
.ends RRE04EA6DFH


******************************************************************************
* Zener Diode
******************************************************************************

.subckt MM3Z4V7ST1G a c
D1 a c zener
C1 a c 200p
.model zener D(BV=4.7)
.ends MM3Z4V7ST1G


******************************************************************************
* Generic DPDT Relay
* Parameter <side> toggles between the A side (0) and B side (1).
******************************************************************************

.subckt DPDT_RELAY coil+ la lc lb rb rc ra coil-
.param side = 0
.param a = !side
.param b = !a

Rlac la lc {a * 100m + b * 10G}
Rrac ra rc {a * 100m + b * 10G}
Clac la lc {a * 100f}
Crac ra rc {a * 100f}

Rlbc lb lc {b * 100m + a * 10G}
Rrbc rb rc {b * 100m + a * 10G}
Clbc lb lc {b * 100f}
Crbc rb rc {b * 100f}
.ends DPDT_RELAY


******************************************************************************
* Generic DPDT Switch
* Parameter <side> toggles between the A side (0) and B side (1).
******************************************************************************

.subckt DPDT_SWITCH a1 c1 b1 a2 c2 b2
.param side = 0
.param a = !side
.param b = !a

Rac1 c1 a1 {a * 100m + b * 10G}
Rac2 c2 a2 {a * 100m + b * 10G}
Cac1 c1 a1 {a * 100f}
Cac2 c2 a2 {a * 100f}

Rbc1 c1 b1 {b * 100m + a * 10G}
Rbc2 c2 b2 {b * 100m + a * 10G}
Cbc1 c1 b1 {b * 100f}
Cbc2 c2 b2 {b * 100f}
.ends DPDT_SWITCH


******************************************************************************
* Digital Potentiometer
******************************************************************************

.subckt DIGIPOT left wiper right
.param value = 25k
.param limit = 100k
.param Cp = 75p
R1 wiper left {value}
C1 wiper left {Cp}
R2 wiper right {limit - value}
C2 wiper right {Cp}
.ends
